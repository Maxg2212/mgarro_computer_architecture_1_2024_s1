package alu_defs;

// Operaciones de la ALU

		parameter ARITH_SUM = 3'b000;
		parameter ARITH_RES = 3'b001;
		parameter ARITH_MUL = 3'b010;
		parameter LOGIC_DLD = 3'b011;
		parameter CR_ = 3'b100;
		
endpackage 